 /*                                                                      
  *  Copyright (c) 2018-2019 Nuclei System Technology, Inc.              
  *  All rights reserved.                                                
  */                                                                     
                                                                         









`ifdef FAKE_FLASH_MODEL
module fake_qspi0_model(
  input  [32-1:2] model_addr, 
  output [32-1:0] model_dout  
  );
        

  wire [31:0] m [0:52-1];




  assign model_dout = m[model_addr[7:2]] 

assign
{
m[00][7:0], m[00][15:8], m[00][23:16], m[00][31:24],
m[01][7:0], m[01][15:8], m[01][23:16], m[01][31:24],
m[02][7:0], m[02][15:8], m[02][23:16], m[02][31:24],
m[03][7:0], m[03][15:8], m[03][23:16], m[03][31:24],
m[04][7:0], m[04][15:8], m[04][23:16], m[04][31:24],
m[05][7:0], m[05][15:8], m[05][23:16], m[05][31:24],
m[06][7:0], m[06][15:8], m[06][23:16], m[06][31:24],
m[07][7:0], m[07][15:8], m[07][23:16], m[07][31:24],
m[08][7:0], m[08][15:8], m[08][23:16], m[08][31:24],
m[09][7:0], m[09][15:8], m[09][23:16], m[09][31:24],

m[10][7:0], m[10][15:8], m[10][23:16], m[10][31:24],
m[11][7:0], m[11][15:8], m[11][23:16], m[11][31:24],
m[12][7:0], m[12][15:8], m[12][23:16], m[12][31:24],
m[13][7:0], m[13][15:8], m[13][23:16], m[13][31:24],
m[14][7:0], m[14][15:8], m[14][23:16], m[14][31:24],
m[15][7:0], m[15][15:8], m[15][23:16], m[15][31:24],
m[16][7:0], m[16][15:8], m[16][23:16], m[16][31:24],
m[17][7:0], m[17][15:8], m[17][23:16], m[17][31:24],
m[18][7:0], m[18][15:8], m[18][23:16], m[18][31:24],
m[19][7:0], m[19][15:8], m[19][23:16], m[19][31:24],

m[20][7:0], m[20][15:8], m[20][23:16], m[20][31:24],
m[21][7:0], m[21][15:8], m[21][23:16], m[21][31:24],
m[22][7:0], m[22][15:8], m[22][23:16], m[22][31:24],
m[23][7:0], m[23][15:8], m[23][23:16], m[23][31:24],
m[24][7:0], m[24][15:8], m[24][23:16], m[24][31:24],
m[25][7:0], m[25][15:8], m[25][23:16], m[25][31:24],
m[26][7:0], m[26][15:8], m[26][23:16], m[26][31:24],
m[27][7:0], m[27][15:8], m[27][23:16], m[27][31:24],
m[28][7:0], m[28][15:8], m[28][23:16], m[28][31:24],
m[29][7:0], m[29][15:8], m[29][23:16], m[29][31:24],

m[30][7:0], m[30][15:8], m[30][23:16], m[30][31:24],
m[31][7:0], m[31][15:8], m[31][23:16], m[31][31:24],
m[32][7:0], m[32][15:8], m[32][23:16], m[32][31:24],
m[33][7:0], m[33][15:8], m[33][23:16], m[33][31:24],
m[34][7:0], m[34][15:8], m[34][23:16], m[34][31:24],
m[35][7:0], m[35][15:8], m[35][23:16], m[35][31:24],
m[36][7:0], m[36][15:8], m[36][23:16], m[36][31:24],
m[37][7:0], m[37][15:8], m[37][23:16], m[37][31:24],
m[38][7:0], m[38][15:8], m[38][23:16], m[38][31:24],
m[39][7:0], m[39][15:8], m[39][23:16], m[39][31:24],

m[40][7:0], m[40][15:8], m[40][23:16], m[40][31:24],
m[41][7:0], m[41][15:8], m[41][23:16], m[41][31:24],
m[42][7:0], m[42][15:8], m[42][23:16], m[42][31:24],
m[43][7:0], m[43][15:8], m[43][23:16], m[43][31:24],
m[44][7:0], m[44][15:8], m[44][23:16], m[44][31:24],
m[45][7:0], m[45][15:8], m[45][23:16], m[45][31:24],
m[46][7:0], m[46][15:8], m[46][23:16], m[46][31:24],
m[47][7:0], m[47][15:8], m[47][23:16], m[47][31:24],
m[48][7:0], m[48][15:8], m[48][23:16], m[48][31:24],
m[49][7:0], m[49][15:8], m[49][23:16], m[49][31:24],

m[50][7:0], m[50][15:8], m[50][23:16], m[50][31:24],
m[51][7:0], m[51][15:8], m[51][23:16], m[51][31:24] 
} =
{
8'h97 ,8'h11 ,8'h00 ,8'h70 ,8'h93 ,8'h81 ,8'h81 ,8'h0A ,8'h17 ,8'h81 ,8'h00 ,8'h70 ,8'h13 ,8'h01 ,8'h81 ,8'hFF,
8'h17 ,8'h05 ,8'h00 ,8'h60 ,8'h13 ,8'h05 ,8'h05 ,8'hFF ,8'h97 ,8'h05 ,8'h00 ,8'h60 ,8'h93 ,8'h85 ,8'h85 ,8'hFE,
8'h63 ,8'h00 ,8'hB5 ,8'h02 ,8'h17 ,8'h16 ,8'h01 ,8'h60 ,8'h13 ,8'h06 ,8'h06 ,8'hFE ,8'h63 ,8'hFA ,8'hC5 ,8'h00,
8'h83 ,8'h22 ,8'h05 ,8'h00 ,8'h23 ,8'hA0 ,8'h55 ,8'h00 ,8'h11 ,8'h05 ,8'h91 ,8'h05 ,8'hE3 ,8'hEA ,8'hC5 ,8'hFE,
8'h17 ,8'h15 ,8'h01 ,8'h60 ,8'h13 ,8'h05 ,8'h45 ,8'hFC ,8'h97 ,8'h05 ,8'h00 ,8'h70 ,8'h93 ,8'h85 ,8'h85 ,8'hFB,
8'h17 ,8'h16 ,8'h00 ,8'h70 ,8'h13 ,8'h06 ,8'h06 ,8'h8D ,8'h63 ,8'hFA ,8'hC5 ,8'h00 ,8'h83 ,8'h22 ,8'h05 ,8'h00,
8'h23 ,8'hA0 ,8'h55 ,8'h00 ,8'h11 ,8'h05 ,8'h91 ,8'h05 ,8'hE3 ,8'hEA ,8'hC5 ,8'hFE ,8'h17 ,8'h15 ,8'h00 ,8'h70,
8'h13 ,8'h05 ,8'h45 ,8'h8B ,8'h97 ,8'h15 ,8'h00 ,8'h70 ,8'h93 ,8'h85 ,8'hC5 ,8'h90 ,8'h63 ,8'h77 ,8'hB5 ,8'h00,
8'h23 ,8'h20 ,8'h05 ,8'h00 ,8'h11 ,8'h05 ,8'hE3 ,8'h6D ,8'hB5 ,8'hFE ,8'h17 ,8'h45 ,8'h00 ,8'h60 ,8'h13 ,8'h05,
8'hA5 ,8'hE1 ,8'h17 ,8'h43 ,8'h00 ,8'h60 ,8'hE7 ,8'h00 ,8'hA3 ,8'hDC ,8'h17 ,8'h43 ,8'h00 ,8'h60 ,8'hE7 ,8'h00,
8'hA3 ,8'hE6 ,8'h99 ,8'h62 ,8'h73 ,8'hA0 ,8'h02 ,8'h30 ,8'h73 ,8'h23 ,8'h00 ,8'h30 ,8'h33 ,8'h73 ,8'h53 ,8'h00,
8'h63 ,8'h02 ,8'h03 ,8'h00 ,8'h01 ,8'h45 ,8'h81 ,8'h45 ,8'h17 ,8'h03 ,8'h00 ,8'h60 ,8'hE7 ,8'h00 ,8'h83 ,8'hF4,
8'h17 ,8'h43 ,8'h00 ,8'h60 ,8'h67 ,8'h00 ,8'h03 ,8'hDB ,8'h01 ,8'hA0 ,8'h00 ,8'h00 ,8'h00 ,8'h00 ,8'h00 ,8'h00  
};

endmodule

`endif
